// $Id: ovm_subscriber.svh,v 1.2 2007/12/14 10:18:56 redelman Exp $
//----------------------------------------------------------------------
//   Copyright 2007-2008 Mentor Graphics Corporation
//   Copyright 2007-2008 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

// This class provides an analysis export. A subclass needs
// to define its own write method Can be useful for
// functional coverage, where the write method will call one
// or more cov.sample methods

// ovm_subscriber - specializations 
// File /usr/local/cds/ovm-2.0/src/methodology/ovm_subscriber.svh, line 27. 
// Original header declaration: 
//   virtual class ovm_subscriber  #( type T = int )



