//----------------------------------------------------------------------
//   Copyright 2007-2008 Mentor Graphics Corporation
//   Copyright 2007-2008 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------


// sequencer_analysis_fifo - specializations 
// File /usr/local/cds/ovm-2.0/src/methodology/sequences/ovm_sequencer_analysis_fifo.svh, line 22. 
// Original header declaration: 
//   class sequencer_analysis_fifo  #(type RSP = ovm_sequence_item)
`include "sequencer_analysis_fifo_ovm_sequence_item.svi"


