// $Id: //dvt/vtech/dev/main/ovm/src/methodology/ovm_pair.svh#5 $
//----------------------------------------------------------------------
//   Copyright 2007-2008 Mentor Graphics Corporation
//   Copyright 2007-2008 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

`ifndef OVM_PAIR_SVH
`define OVM_PAIR_SVH

//
// paramterized pair classes
//

// ovm_class_pair - specializations 
// File /usr/local/cds/ovm-2.0/src/methodology/ovm_pair.svh, line 29. 
// Original header declaration: 
//   class ovm_class_pair  #( type T1 = int ,
// 			type T2 = T1 )



// ovm_built_in_pair - specializations 
// File /usr/local/cds/ovm-2.0/src/methodology/ovm_pair.svh, line 95. 
// Original header declaration: 
//   class ovm_built_in_pair  #( type T1 = int ,
// 			   type T2 = T1 )



`endif // OVM_PAIR_SVH
