module overlapController(clk);
	
	parameter halfWindowSize = 512;
	parameter wordLength = 16;
	
	input clk;
	
	
	always @(posedge clk )
	begin 
	
	end
	
endmodule
