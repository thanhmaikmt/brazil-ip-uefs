// $Id: ovm_ports.svh,v 1.7 2008/07/18 10:15:20 redelman Exp $
//----------------------------------------------------------------------
//   Copyright 2007-2008 Mentor Graphics Corporation
//   Copyright 2007-2008 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

// ovm_blocking_put_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 22. 
// Original header declaration: 
//   class ovm_blocking_put_port  #(type T=int)

 

// ovm_nonblocking_put_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 28. 
// Original header declaration: 
//   class ovm_nonblocking_put_port  #(type T=int)



// ovm_put_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 34. 
// Original header declaration: 
//   class ovm_put_port  #(type T=int)
`include "ovm_put_port_stream.svi"
`include "ovm_put_port_amostra.svi"
`include "ovm_put_port_erro.svi"



// ovm_blocking_get_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 40. 
// Original header declaration: 
//   class ovm_blocking_get_port  #(type T=int)

 

// ovm_nonblocking_get_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 46. 
// Original header declaration: 
//   class ovm_nonblocking_get_port  #(type T=int)



// ovm_get_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 52. 
// Original header declaration: 
//   class ovm_get_port  #(type T=int)
`include "ovm_get_port_stream.svi"
`include "ovm_get_port_amostra.svi"
`include "ovm_get_port_erro.svi"

 

// ovm_blocking_peek_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 58. 
// Original header declaration: 
//   class ovm_blocking_peek_port  #(type T=int)

 

// ovm_nonblocking_peek_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 64. 
// Original header declaration: 
//   class ovm_nonblocking_peek_port  #(type T=int)



// ovm_peek_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 70. 
// Original header declaration: 
//   class ovm_peek_port  #(type T=int)

 

// ovm_blocking_get_peek_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 76. 
// Original header declaration: 
//   class ovm_blocking_get_peek_port  #(type T=int)

 

// ovm_nonblocking_get_peek_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 82. 
// Original header declaration: 
//   class ovm_nonblocking_get_peek_port  #(type T=int)



// ovm_get_peek_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 88. 
// Original header declaration: 
//   class ovm_get_peek_port  #(type T=int)

 

// ovm_blocking_master_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 94. 
// Original header declaration: 
//   class ovm_blocking_master_port  #(type REQ=int, type RSP=int)

 

// ovm_nonblocking_master_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 101. 
// Original header declaration: 
//   class ovm_nonblocking_master_port  #(type REQ=int, type RSP=int)

 

// ovm_master_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 108. 
// Original header declaration: 
//   class ovm_master_port  #(type REQ=int, type RSP=int)



// ovm_blocking_slave_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 115. 
// Original header declaration: 
//   class ovm_blocking_slave_port  #(type REQ=int, type RSP=int)

 

// ovm_nonblocking_slave_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 122. 
// Original header declaration: 
//   class ovm_nonblocking_slave_port  #(type REQ=int, type RSP=int)

 

// ovm_slave_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 129. 
// Original header declaration: 
//   class ovm_slave_port  #(type REQ=int, type RSP=int)



// ovm_blocking_transport_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 136. 
// Original header declaration: 
//   class ovm_blocking_transport_port  #(type REQ=int, type RSP=int)



// ovm_nonblocking_transport_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 142. 
// Original header declaration: 
//   class ovm_nonblocking_transport_port  #(type REQ=int, type RSP=int)



// ovm_transport_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 148. 
// Original header declaration: 
//   class ovm_transport_port  #(type REQ=int, type RSP=int)



// ovm_analysis_port - specializations 
// File /usr/local/cds/ovm-2.0/src/tlm/ovm_ports.svh, line 154. 
// Original header declaration: 
//   class ovm_analysis_port  # (type T = int)
`include "ovm_analysis_port_ovm_sequence_item.svi"
`include "ovm_analysis_port_stream.svi"
`include "ovm_analysis_port_amostra.svi"
`include "ovm_analysis_port_erro.svi"


