// $Id: //dvt/vtech/dev/main/ovm/src/base/ovm_registry.svh#14 $
//----------------------------------------------------------------------
//   Copyright 2007-2008 Mentor Graphics Corporation
//   Copyright 2007-2008 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------
`ifndef OVM_REGISTRY_SVH
`define OVM_REGISTRY_SVH

// ovm_component_registry - specializations 
// File /usr/local/cds/ovm-2.0/src/base/ovm_registry.svh, line 24. 
// Original header declaration: 
//   class ovm_component_registry  #(type T=ovm_component, string Tname="<unknown>")




// ovm_object_registry - specializations 
// File /usr/local/cds/ovm-2.0/src/base/ovm_registry.svh, line 82. 
// Original header declaration: 
//   class ovm_object_registry  #(type T=ovm_object, string Tname="<unknown>")



`endif
