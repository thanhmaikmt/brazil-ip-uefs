// $Id: ovm_random_stimulus.svh,v 1.5 2008/08/19 10:13:23 redelman Exp $
//----------------------------------------------------------------------
//   Copyright 2007-2008 Mentor Graphics Corporation
//   Copyright 2007-2008 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------


// A general purpose unidirectional random stimulus class.
//
// If you want to do stuff before or after the run method,
// extend this class, define your own run, and call
// super.run( . ). This will be the case, for example when
// you need a non random initialisation sequence before you
// do some constraint random testing.
//

// The ovm_stimulus class generates streams of trans_type
// transactions. These streams may be generated by the
// randomize method of trans_type, or the randomize method
// of one of its subclasses.  The stream may go
// indefinitely, until terminated by a call to
// stop_stimulus_generation, or we may specify the maximum
// number of transactions to be generated.
//
// By using inheritance, we can add directed initialization
// or tidy up sequences to the random stimulus generation.

// ovm_random_stimulus - specializations 
// File /usr/local/cds/ovm-2.0/src/methodology/ovm_random_stimulus.svh, line 43. 
// Original header declaration: 
//   class ovm_random_stimulus  #(type trans_type=ovm_transaction)


