// $Id: ovm_scenario_driver.svh,v 1.9 2008/08/07 15:18:05 jlrose Exp $
//----------------------------------------------------------------------
//   Copyright 2007-2008 Mentor Graphics Corporation
//   Copyright 2007-2008 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------


//typedef class ovm_scenario_controller_base;
//typedef class ovm_scenario_base;

// ovm_scenario_driver - specializations 
// File /usr/local/cds/ovm-2.0/src/methodology/layered_stimulus/ovm_scenario_driver.svh, line 26. 
// Original header declaration: 
//   virtual class ovm_scenario_driver  #(type REQ = ovm_sequence_item, type RSP = REQ)



